//
// Copyright (c) 2015-2016 Jong Hun Han
// Copyright (c) 2015 SRI International
// All rights reserved
//
// This software was developed by Stanford University and the University of
// Cambridge Computer Laboratory under National Science Foundation under Grant
// No. CNS-0855268, the University of Cambridge Computer Laboratory under EPSRC
// INTERNET Project EP/H040536/1 and by the University of Cambridge Computer
// Laboratory under DARPA/AFRL contract FA8750-11-C-0249 ("MRC2"), as part of
// the DARPA MRC research programme.
//
// @NETFPGA_LICENSE_HEADER_START@
//
// Licensed to NetFPGA C.I.C. (NetFPGA) under one or more contributor license
// agreements.  See the NOTICE file distributed with this work for additional
// information regarding copyright ownership.  NetFPGA licenses this file to you
// under the NetFPGA Hardware-Software License, Version 1.0 (the "License"); you
// may not use this file except in compliance with the License.  You may obtain
// a copy of the License at:
//
//   http://www.netfpga-cic.org
//
// Unless required by applicable law or agreed to in writing, Work distributed
// under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied.  See the License for the
// specific language governing permissions and limitations under the License.
//
// @NETFPGA_LICENSE_HEADER_END@

`timescale 1ns/1ps

`include "nf_sume_blueswitch_register_define.v"
`include "nf_sume_blueswitch_parameter_define.v"

module tcam_multi_wrapper
#(
   parameter   TCAM_ADDR_WIDTH   = 5,
   parameter   TCAM_DATA_WIDTH   = 32
)
(
   input                                     CLK,
   input                                     RSTN,

   input                                     WR,
   input          [TCAM_ADDR_WIDTH-1:0]      ADDR_WR,
   input          [TCAM_DATA_WIDTH-1:0]      DIN,
   input          [TCAM_DATA_WIDTH-1:0]      DIN_MASK,
   output   wire                             BUSY,

`ifdef EN_TCAM_RD
   input                                     RD,
   input          [TCAM_ADDR_WIDTH-1:0]      ADDR_RD,
   output   reg   [TCAM_DATA_WIDTH-1:0]      DOUT,
`endif

   input          [TCAM_DATA_WIDTH-1:0]      CAM_DIN,
   input          [TCAM_DATA_WIDTH-1:0]      CAM_DATA_MASK,
   output   wire                             MATCH,
   output   wire  [TCAM_ADDR_WIDTH-1:0]      MATCH_ADDR
);

`ifdef XIL_TCAM_USE
//Use TCAM macro blocks generated by Xilinx tool.
//

reg   [TCAM_ADDR_WIDTH-2:0]   rADDR_WR_0, rADDR_WR_1;
reg   [TCAM_DATA_WIDTH-1:0]   rDIN, rDIN_MASK, rCAM_DIN, rCAM_DATA_MASK;
reg   rWR_0, rWR_1;
`ifdef EN_TCAM_RD
reg   rRD;
reg   [TCAM_ADDR_WIDTH-2:0]   rADDR_RD;
`endif

always @(posedge CLK)
   if (~RSTN) begin
      rWR_0             <= 0;
      rWR_1             <= 0;
      `ifdef EN_TCAM_RD
      rRD               <= 0;
      rADDR_RD          <= 0;
      `endif
      rADDR_WR_0        <= 0;
      rADDR_WR_1        <= 0;
      rDIN              <= 0;
      rDIN_MASK         <= 0;
      rCAM_DIN          <= 0;
      rCAM_DATA_MASK    <= 0;
   end
   else begin
      rWR_0             <= WR & ~ADDR_WR[TCAM_ADDR_WIDTH-1];
      rWR_1             <= WR & ADDR_WR[TCAM_ADDR_WIDTH-1];
      `ifdef EN_TCAM_RD
      rRD               <= RD;
      rADDR_RD          <= ADDR_RD;
      `endif
      rADDR_WR_0        <= ADDR_WR[TCAM_ADDR_WIDTH-2:0];
      rADDR_WR_1        <= ADDR_WR[TCAM_ADDR_WIDTH-2:0];
      rDIN              <= DIN;
      rDIN_MASK         <= DIN_MASK;
      rCAM_DIN          <= CAM_DIN;
      rCAM_DATA_MASK    <= CAM_DATA_MASK;
   end

wire  [TCAM_ADDR_WIDTH-2:0]   wMATCH_ADDR_0, wMATCH_ADDR_1;
wire  wMATCH_0, wMATCH_1, wBUSY_0, wBUSY_1;

reg   [TCAM_ADDR_WIDTH-2:0]   rMATCH_ADDR_0, rMATCH_ADDR_1;
reg   rMATCH_0, rMATCH_1, rBUSY_0, rBUSY_1;

always @(posedge CLK)
   if (~RSTN) begin
      rBUSY_0        <= 0;
      rMATCH_0       <= 0;
      rMATCH_ADDR_0  <= 0;
      rBUSY_1        <= 0;
      rMATCH_1       <= 0;
      rMATCH_ADDR_1  <= 0;
  end
   else begin
      rBUSY_0        <= wBUSY_0;
      rMATCH_0       <= wMATCH_0;
      rMATCH_ADDR_0  <= wMATCH_ADDR_0;
      rBUSY_1        <= wBUSY_1;
      rMATCH_1       <= wMATCH_1;
      rMATCH_ADDR_1  <= wMATCH_ADDR_1;
   end

assign BUSY = rBUSY_0 | rBUSY_1;
assign MATCH = rMATCH_0 | rMATCH_1;
assign MATCH_ADDR = (rMATCH_0) ? {1'b0, rMATCH_ADDR_0} : (rMATCH_1) ? {1'b1, rMATCH_ADDR_1} : 0;


nf_sume_tcam
#(
   .C_TCAM_ADDR_WIDTH   (  TCAM_ADDR_WIDTH-1 ),
   .C_TCAM_DATA_WIDTH   (  TCAM_DATA_WIDTH   )
)
tcam_0
(
   .CLK                 (  CLK               ), 
   .DIN                 (  rDIN              ), 
   .WE                  (  rWR_0             ), 
   .WR_ADDR             (  rADDR_WR_0        ),

   .BUSY                (  wBUSY_0           ), 
   .MATCH               (  wMATCH_0          ), 
   .MATCH_ADDR          (  wMATCH_ADDR_0     ),
   .DATA_MASK           (  {(TCAM_DATA_WIDTH){1'b1}} ), 
   //.DATA_MASK           (  rDIN_MASK         ), 
   .CMP_DIN             (  rCAM_DIN          ),
   .CMP_DATA_MASK       (  rCAM_DATA_MASK    )
   //.CMP_DATA_MASK       (  {(TCAM_DATA_WIDTH){1'b1}} )
);

nf_sume_tcam
#(
   .C_TCAM_ADDR_WIDTH   (  TCAM_ADDR_WIDTH-1 ),
   .C_TCAM_DATA_WIDTH   (  TCAM_DATA_WIDTH   )
)
tcam_1
(
   .CLK                 (  CLK               ), 
   .DIN                 (  rDIN              ), 
   .WE                  (  rWR_1             ), 
   .WR_ADDR             (  rADDR_WR_1        ),

   .BUSY                (  wBUSY_1           ), 
   .MATCH               (  wMATCH_1          ), 
   .MATCH_ADDR          (  wMATCH_ADDR_1     ),
   .DATA_MASK           (  {(TCAM_DATA_WIDTH){1'b1}} ), 
   //.DATA_MASK           (  rDIN_MASK         ), 
   .CMP_DIN             (  rCAM_DIN          ),
   .CMP_DATA_MASK       (  rCAM_DATA_MASK    )
   //.CMP_DATA_MASK       (  {(TCAM_DATA_WIDTH){1'b1}} )
);

//generate
//   if (TCAM_ADDR_WIDTH == 5) begin
//      if (TCAM_DATA_WIDTH == 16) begin : tcam_16x16
//         tcam16x16 tcam16x16_0 (
//            .CLK           (  CLK               ), 
//            .WE            (  rWR_0             ), 
//            .BUSY          (  wBUSY_0           ), 
//            .MATCH         (  wMATCH_0          ), 
//            .DIN           (  rDIN              ), 
//            .DATA_MASK     (  rDIN_MASK         ), 
//            .WR_ADDR       (  rADDR_WR_0        ),
//            .CMP_DIN       (  rCAM_DIN          ),
//            .CMP_DATA_MASK (  rCAM_DATA_MASK    ),
//            .MATCH_ADDR    (  wMATCH_ADDR_0     )
//         );
//
//         tcam16x16 tcam16x16_1 (
//            .CLK           (  CLK               ), 
//            .WE            (  rWR_1             ), 
//            .BUSY          (  wBUSY_1           ), 
//            .MATCH         (  wMATCH_1          ), 
//            .DIN           (  rDIN              ), 
//            .DATA_MASK     (  rDIN_MASK         ), 
//            .WR_ADDR       (  rADDR_WR_1        ),
//            .CMP_DIN       (  rCAM_DIN          ),
//            .CMP_DATA_MASK (  rCAM_DATA_MASK    ),
//            .MATCH_ADDR    (  wMATCH_ADDR_1     )
//         );
//      end
//      else if (TCAM_DATA_WIDTH == 32) begin : tcam_16x32
//         tcam16x32 tcam16x32_0 (
//            .CLK           (  CLK               ), 
//            .WE            (  rWR_0             ), 
//            .BUSY          (  wBUSY_0           ), 
//            .MATCH         (  wMATCH_0          ), 
//            .DIN           (  rDIN              ), 
//            .DATA_MASK     (  rDIN_MASK         ), 
//            .WR_ADDR       (  rADDR_WR_0        ),
//            .CMP_DIN       (  rCAM_DIN          ),
//            .CMP_DATA_MASK (  rCAM_DATA_MASK    ),
//            .MATCH_ADDR    (  wMATCH_ADDR_0     )
//         );
//
//         tcam16x32 tcam16x32_1 (
//            .CLK           (  CLK               ), 
//            .WE            (  rWR_1             ), 
//            .BUSY          (  wBUSY_1           ), 
//            .MATCH         (  wMATCH_1          ), 
//            .DIN           (  rDIN              ), 
//            .DATA_MASK     (  rDIN_MASK         ), 
//            .WR_ADDR       (  rADDR_WR_1        ),
//            .CMP_DIN       (  rCAM_DIN          ),
//            .CMP_DATA_MASK (  rCAM_DATA_MASK    ),
//            .MATCH_ADDR    (  wMATCH_ADDR_1     )
//         );
//      end
//      else if (TCAM_DATA_WIDTH == 48) begin : tcam_16x48
//         tcam16x48 tcam16x48_0 (
//            .CLK           (  CLK               ), 
//            .WE            (  rWR_0             ), 
//            .BUSY          (  wBUSY_0           ), 
//            .MATCH         (  wMATCH_0          ), 
//            .DIN           (  rDIN              ), 
//            .DATA_MASK     (  rDIN_MASK         ), 
//            .WR_ADDR       (  rADDR_WR_0        ),
//            .CMP_DIN       (  rCAM_DIN          ),
//            .CMP_DATA_MASK (  rCAM_DATA_MASK    ),
//            .MATCH_ADDR    (  wMATCH_ADDR_0     )
//         );
//
//         tcam16x48 tcam16x48_1 (
//            .CLK           (  CLK               ), 
//            .WE            (  rWR_1             ), 
//            .BUSY          (  wBUSY_1           ), 
//            .MATCH         (  wMATCH_1          ), 
//            .DIN           (  rDIN              ), 
//            .DATA_MASK     (  rDIN_MASK         ), 
//            .WR_ADDR       (  rADDR_WR_1        ),
//            .CMP_DIN       (  rCAM_DIN          ),
//            .CMP_DATA_MASK (  rCAM_DATA_MASK    ),
//            .MATCH_ADDR    (  wMATCH_ADDR_1     )
//         );
//      end
//   end
//endgenerate

`else
//This is simple register based TCAM design, which is not recommneded
//due to increasing costs of fpga resources.

reg   [TCAM_ADDR_WIDTH-1:0]   rADDR_WR, rMATCH_ADDR;
reg   [TCAM_DATA_WIDTH-1:0]   rDIN;
reg   [TCAM_DATA_WIDTH-1:0]   rCAM_DIN;
reg   rWR, rBUSY, rMATCH;

wire  [TCAM_ADDR_WIDTH-1:0]   wMATCH_ADDR;
wire  wMATCH;

assign BUSY = rBUSY;
assign MATCH = rMATCH;
assign MATCH_ADDR = rMATCH_ADDR;

always @(posedge CLK)
   if (~RSTN) begin
      rWR         <= 0;
      rADDR_WR    <= 0;
      rDIN        <= 0;
      rCAM_DIN    <= 0;
   end
   else begin
      rWR         <= WR;
      rADDR_WR    <= ADDR_WR;
      rDIN        <= DIN;
      rCAM_DIN    <= CAM_DIN;
   end

always @(posedge CLK)
   if (~RSTN) begin
      rBUSY       <= 0;
      rMATCH      <= 0;
      rMATCH_ADDR <= 0;
   end
   else begin
      rBUSY       <= WR | rWR;
      rMATCH      <= wMATCH;
      rMATCH_ADDR <= wMATCH_ADDR;
   end


tcam_rtl
#(
   .ADDR_WIDTH    (  TCAM_ADDR_WIDTH         ),
   .DATA_WIDTH    (  TCAM_DATA_WIDTH         )
)
tcam_rtl
(
   .CLK           (  CLK                     ),
   .WR            (  rWR                     ),
   .ADDR_WR       (  rADDR_WR                ),
   .DIN           (  rDIN                    ),
   .DIN_MASK      (  {TCAM_DATA_WIDTH{1'b1}} ),

`ifdef EN_TCAM_RD
   .RD            (  0                       ),
   .ADDR_RD       (  0                       ),
   .DOUT          (                          ),
`endif

   .CAM_IN        (  rCAM_DIN                ),
   .MATCH         (  wMATCH                  ),
   .MATCH_ADDR    (  wMATCH_ADDR             )
);

`endif


endmodule
